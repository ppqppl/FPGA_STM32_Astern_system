module beep_driver (
    input   wire          clk     ,
    input   wire          rstn    ,

    output  wire          beep    
);



endmodule //beep_driver